`default_nettype none
`timescale 1ns / 1ps

module hybrid_synthesis_tb;

logic clk;
logic rst;
logic window_switching_flag_in;
logic [1:0] block_type_in;
logic mixed_block_flag_in;
logic new_frame_start;

logic [31:0] x_in;
logic din_valid;
logic [31:0] x_out;
logic dout_valid;


logic [576 * 32 - 1 :0] CODE;


hybrid_synthesis UUT (
    .clk(clk),
    .rst(rst),
    .window_switching_flag_in(window_switching_flag_in),
    .block_type_in(block_type_in),
    .mixed_block_flag_in(mixed_block_flag_in),
    .new_frame_start(new_frame_start),
    .x_in(x_in),
    .din_valid(din_valid),
    .x_out(x_out),
    .dout_valid(dout_valid)
  );


always begin
  #10;
  clk = !clk;     //clock cycles now happend every 20!
end


initial begin
  $dumpfile("sim/hybrid_synthesis_tb.vcd");
  $dumpvars(0, hybrid_synthesis_tb);
  $display("Starting Sim");

  CODE = 18432'h001879cd000e411f00000000fff1bee1ffdc14cbffcfa274ffc2532cffc2532cffc2532cffc2532cffcfb00affdc4989ffe7c6c8fff25832fffb7773fffc669c0001bc8200027bad000f222a000f3cb9000725070006976e0006fac60006a79f000ec350000e6ee8000e411f000e411f000e4e98000e7491000ed38c00108159000a03d2000d0ac400068ee100027bad000f222a00183ff60015785e001709d10017049b000da891000e0cf0000e3398000e411f0005a82700059aa4ffffcc30ffffc4adffff770b00000000fffc669cfffdae3e00027bad000f222a0007a80a0007250700000000fffa5e56fffa5910fff1bf40fff1b98cfff1bee1fff1bee1fff1cc68fff1f310fff2576ffffbb773fffd07d5ffff18580001bc8200027bad000f222a000f3cb9000f4f21000f0bac000eb9b9000ed38c000e7491000e4e980005a8270005a8270005a8240005a8020005a6f0000518b40004888d00039964000251c20001f0b6fff83d26fff857f6fff8daf9fff96892fff9d561ffffc4adffffeb71fffffaa5000000000000000000000000ffffeb7100056b9d0004488d00011c290005ddc0000105cdffffa15effe3adaaffe3b1c6ffe44a44ffe6e74ffff14647fffa1dbdfffa57fe000000000005a827000e411f000e4e98000e7491000ed38c000f89e0000827d00009d6c20006b96800027bad000f222a000c9195000bc37e000cfccc000cd7a7000da891000e0cf0000e3398000e411f000e411f000e4674000e5550000e7962000eb9b90006976e000725070002ab240002e9110004d9c80004fce6000399640004888d0004488d000511730005743100059aa40005a8270005a8270000000000000000000000000000000000000000fffaa0cbfffb031a0002e9110004d9c80002ab240001c5d100000000000000000000000000000000000000000000000000000000000000000000000000003b53000088f5000107700001c5d10002ab24fffe0f4a0007c2da0004fce600055f3500058ffe0005a1aa0005a6f0000000000000000000000000fffa57d9fffa5d37fffa6c8efffa9463fffae74cfffb7773fffc669cfffdae3efffe0f4a0007c2da0007a80a000725070006976e00062a9f0005e2430005bc920005ad800005a8270000000000000000ffffeb71ffffc4adffff770bfffef890fffe3a2f000251c2fffd16effffb2638fff857f6fffaa0cbfffa7002fffa5e56fffa5910fffa57fe0000000000000000000000000000055b0005bc920005e24300062a9f0006976e0001c5d10002ab240002e9110004d9c80004fce600055f350004888d000518b400056b9d000593720005a8240005a8270005a8270005a2c90005937200056b9d000518b40004888d00039964000251c20001f0b6fff83d26fff857f6fff8daf9fff96892fff9d561fffa1dbdfffa436efffa5280fffa57d9fffa57d9fffa5d37fffa6c8efffa9463fffae74cfffb7773fffc669cfffdae3efffe0f4a0007c2da0007a80a000725070006976e00062a9f0005e2430005bc920005ad800000000000000000fffffaa5ffffeb71ffffc4ad00000000000000000000000000000000000000000000000000000000000000000000000000000000fffa5910fffa57fefffa57dcfffa57d9fffa57d9fffa57dcfffa57fefffa5910fffa5e5600000000000000000002ab240002e9110004d9c80004fce60000000000000000000088f500003b530000148f0000055b0000000000000000000000000000000000000000000000000000000000000000fffd54dcfffd16effffb2638fffb031a000000000000000000000000000000000000000000000000000000000005a8270005ad800005bc920005e2430000000000000000000000000000000000000000000000000000000000000000000000000000000000056b9d000593720005a2c90005a8270005a8270005a2c90005937200056b9d000518b40004888d00039964000251c20001f0b6fff83d26fff857f6fff8daf9fff96892fff9d561fffa1dbdfffa436efffa5280000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000107700001c5d10002ab240002e9110004d9c80004fce600055f3500058ffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;



  clk = 0;
  rst = 0;
  x_in = 0;
  window_switching_flag_in = 1;
  block_type_in = 1;
  mixed_block_flag_in = 0;
  new_frame_start = 0;
  din_valid = 0;
  #20;
  rst = 1;
  #20;
  rst = 0;
  #20

  din_valid = 1;
  for (int i = 0; i < 576; i ++) begin
    x_in = CODE >> ((576 - 1 - i) * 32);
    #20;
  end

  CODE = 18432'h14d4471403649d14edf8291d04d065f8fde420ccfcd4ce55fe16ec20fcd4ce55fc9b62ecff9a6806ff9a68060088cc4e00bb0a3c0095c41b007a44f800c7efe7001428a200d92745ff9e18cc0095c41bfefa5d3fffae106bff3c4a2dffb51df3ffbb99d9fffa57d9ff80000100446627ff86207500229d2e0032cbfdffb4407600229d2eff3c4a2dff86207500446627ffd7aebbfff4afb1ffbac5a400ae718eff9f44e7fea74a5d00d63f8f001c823d000fffffffbac5a4007b59a900ae718efff0000100977f1400977f1400000000007b59a9000b504f00453a5c0030f39a0114c6adfea74a5d0060bb190047d66affd7aebb00000000ffe37dc3006597fa001c823dff9f44e7ffcf0c66fff4afb1ffcf0c66ffcf0c660060bb190047d66affcf0c66ffe37dc3ffe37dc3fff4afb1001c823d0030f39a007b59a9000b504f001c823dfff4afb100000000ff84a657000b504f000000000030f39affcf0c660060bb19fff4afb1ffbac5a40047d66affcd340300453a5c0030f39a006b1fc7ffd7aebb0030f39a0032cbfd00285145ff6880ecfff80001ffd7aebbfff4afb1ffebd75e00453a5cfff4afb1ffebd75efff00001ffe37dc3ffdd62d2006597fa001c823dfff80001ff7733b2ffcf0c66ffcd340300453a5cffe37dc3ffebd75e0047d66a0030f39affe37dc3ff6880ec000b504f001c823dff6880ecffb829960030f39a0060bb19ffe37dc30030f39a0047d66a00000000000b504f001c823d001c823d0030f39a0030f39a001c823dffb82996ff9f44e7ffcf0c66ffcf0c66ffe37dc3ffb82996000b504f000b504f0000000000000000001c823dffe37dc3fff4afb1ffb82996001c823d001c823d000fffffffd7aebbffbac5a4000fffff000000000028514500000000fff00001000fffffffd7aebb0028514500285145000fffffffd7aebb000fffff00453a5c000fffff00285145000fffff00453a5cffbac5a400000000ffd7aebb00000000ff9a680600453a5cffd7aebbff9a6806ffbac5a4ffd7aebb00453a5c00000000fff00001fff00001fff00001fff00001006597faffbac5a4006597fa00453a5c00285145ffbac5a4000fffff00453a5c0060bb19ffd7aebb006597faffcf0c66fff00001ffbac5a4ffb829960000000000285145001c823d00285145fff00001ffcf0c66000fffff000000000000000000453a5c00000000ffcf0c66fff00001000fffffffe37dc3ffbac5a400285145ffe37dc30028514500285145001c823dfff0000100000000ffe37dc3ffbac5a400000000000b504fffd7aebbfff0000100000000000fffff000fffff00000000fff00001ffd7aebb0030f39a000fffff00453a5c001c823dfff0000100000000001c823dfff00001000fffff0000000000285145000b504f00000000ffd7aebbfff4afb1000fffffffbac5a40030f39afff00001fff00001ffcf0c66ffd7aebb00285145000b504f0000000000285145001c823d006597fa000fffff001c823dfff00001000fffff001c823dfff0000100453a5c0000000000000000000fffff000b504ffff0000100000000fff4afb1000fffff000000000030f39afff00001000000000000000000000000000000000047d66a000fffff00000000001c823d000ffffffff000010000000000285145ffd7aebb001c823dffd7aebb00000000fff4afb1fff0000100000000000b504f00000000ffd7aebbfff4afb100000000000000000000000000000000fff00001ffe37dc3000ffffffff4afb1fff4afb1ffebd75efff4afb1000000000007ffff000000000000000000000000001c823d00000000001428a2fff4afb1000b504f00000000001c823dfff4afb1fff80001001c823d00000000fff80001ffe37dc3fff4afb1ffebd75e000b504f00000000001428a2000b504f000b504f00000000ffe37dc3000b504f00000000fff4afb1000b504f001428a200000000001c823d001428a200000000fff4afb100000000000b504f000000000007ffff001c823d000b504f00000000fff4afb1000000000007ffff000b504ffff4afb1000000000000000000000000ffebd75e000b504f000b504f00000000001c823d000b504f00000000fff4afb10000000000000000001c823d000b504ffff800010000000000000000fff800010000000000000000fff8000100000000000b504fffebd75e000b504f000b504f0007ffff00000000fff4afb100000000001c823dfff4afb1ffebd75e00000000000000000007ffff000000000000000000000000fff0000100000000fff00001000ffffffff0000100000000fff0000100000000000fffff00000000fff00001000fffff00000000fff00001000fffff00000000fff0000100000000fff000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

  block_type_in = 2;
  window_switching_flag_in = 1;
  mixed_block_flag_in = 0;

  for (int i = 0; i < 576; i ++) begin
    x_in = CODE >> ((576 - 1 - i) * 32);
    #20;
  end

  din_valid = 0;
  #2000;

  new_frame_start = 1;
  #20;
  new_frame_start = 0;
  #500;

  $display("Finishing Sim");
  $finish;

end
endmodule

`default_nettype wire
