`default_nettype none
`timescale 1ns / 1ps


module HT_30(
		input wire clk,
		input wire rst,
		
		input wire axiiv,
		input wire axiid,
		output logic axiov,
		output logic signed [15:0] x_val,
		output logic signed [15:0] y_val
	);

  parameter MAX_BITS = 12;
	parameter LINBITS =11;

	logic [11:0] buffer;
	logic [4:0] bit_counter;
	logic [3:0] x_linbit_counter, y_linbit_counter;
	logic x_signbit_counter, y_signbit_counter;

	logic [8:0] word;
	logic found;
	logic [3:0] x_abs, y_abs;
	logic x_sign, y_sign;
	logic [LINBITS - 1:0] x_linval, y_linval;

	assign {found, x_abs, y_abs} = word;

	logic [MAX_BITS-2:0] buffer_clearer_with_input;
	assign buffer_clearer_with_input = 0;


	always_comb begin
		x_val = (~x_sign) ? x_abs + x_linval : -8'sd1 * (x_abs + x_linval);
		y_val = (~y_sign) ? y_abs + y_linval : -8'sd1 * (y_abs + y_linval);

		axiov = ( found )
				&& ( (x_abs < 4'd15) || (x_linbit_counter == LINBITS) )
				&& ( (x_abs == 0) || (x_signbit_counter) )
				&& ( (y_abs < 4'd15) || (y_linbit_counter == LINBITS) )
				&& ( (y_abs == 0) || (y_signbit_counter));
	end
	always_ff @(posedge clk) begin
		if (rst) begin
			bit_counter <= 0;
			buffer <= 0;
      x_sign <= 0;
      y_sign <= 0;
      x_linval <= 0;
      y_linval <= 0;
      x_linbit_counter <= 0;
      y_linbit_counter <= 0;
      x_signbit_counter <= 0;
      y_signbit_counter <= 0;
		end else begin
			if (axiov) begin
				bit_counter <= axiiv ? 1 : 0;
				buffer <= axiiv ? {axiid, buffer_clearer_with_input} : 0;
        x_sign <= 0;
        y_sign <= 0;
        x_linval <= 0;
        y_linval <= 0;
        x_linbit_counter <= 0;
        y_linbit_counter <= 0;
        x_signbit_counter <= 0;
        y_signbit_counter <= 0;
      end else if (axiiv) begin
        if (~found) begin
  		    bit_counter <= bit_counter + 1;
  		    case (bit_counter)
						5'd0 : buffer[11] <= axiid;
						5'd1 : buffer[10] <= axiid;
						5'd2 : buffer[9] <= axiid;
						5'd3 : buffer[8] <= axiid;
						5'd4 : buffer[7] <= axiid;
						5'd5 : buffer[6] <= axiid;
						5'd6 : buffer[5] <= axiid;
						5'd7 : buffer[4] <= axiid;
						5'd8 : buffer[3] <= axiid;
						5'd9 : buffer[2] <= axiid;
						5'd10 : buffer[1] <= axiid;
						5'd11 : buffer[0] <= axiid;
          endcase
			
        end else if ((x_abs == 4'd15) && (x_linbit_counter < LINBITS)) begin
          x_linval <= {x_linval[LINBITS - 2:0], axiid};
          x_linbit_counter <= x_linbit_counter + 1;
        end else if ((x_abs > 0) && ~x_signbit_counter) begin
          x_sign <= axiid;
          x_signbit_counter <= x_signbit_counter + 1;
        end else if ((y_abs == 4'd15) && (y_linbit_counter < LINBITS)) begin
          y_linval <= {y_linval[LINBITS - 2:0], axiid};
          y_linbit_counter <= y_linbit_counter + 1;
        end else if ((y_abs > 0) && ~y_signbit_counter) begin
          y_sign <= axiid;
          y_signbit_counter <= y_signbit_counter + 1;
        end
			end
		end
	end
	always_comb begin
		case (bit_counter)
			5'd0 : word = 9'b0_0000_0000;
			5'd1 : word = 10'b00_0000_0000;
			5'd2 : word = 10'b00_0000_0000;
			5'd3 : word = 10'b00_0000_0000;
			5'd4 : begin
					case (buffer[11:8])
						4'b1111 : word = 9'b1_0000_0000;
						4'b1101 : word = 9'b1_0000_0001;
						4'b1110 : word = 9'b1_0001_0000;
						4'b1100 : word = 9'b1_0001_0001;
						4'b0011 : word = 9'b1_1111_1111;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd5 : begin
					case (buffer[11:7])
						5'b10101 : word = 9'b1_0001_0010;
						5'b10110 : word = 9'b1_0010_0001;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd6 : begin
					case (buffer[11:6])
						6'b101110 : word = 9'b1_0000_0010;
						6'b100110 : word = 9'b1_0001_0011;
						6'b101111 : word = 9'b1_0010_0000;
						6'b101001 : word = 9'b1_0010_0010;
						6'b100111 : word = 9'b1_0011_0001;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd7 : begin
					case (buffer[11:5])
						7'b1010000 : word = 9'b1_0000_0011;
						7'b1000111 : word = 9'b1_0001_0100;
						7'b1001010 : word = 9'b1_0010_0011;
						7'b1000100 : word = 9'b1_0010_0100;
						7'b0010010 : word = 9'b1_0010_1111;
						7'b1010001 : word = 9'b1_0011_0000;
						7'b1001011 : word = 9'b1_0011_0010;
						7'b1000110 : word = 9'b1_0011_0011;
						7'b0010000 : word = 9'b1_0011_1111;
						7'b1001000 : word = 9'b1_0100_0001;
						7'b1000101 : word = 9'b1_0100_0010;
						7'b0001110 : word = 9'b1_0100_1111;
						7'b1000010 : word = 9'b1_0101_0001;
						7'b0001100 : word = 9'b1_0101_1111;
						7'b0001010 : word = 9'b1_0110_1111;
						7'b0010100 : word = 9'b1_1111_0001;
						7'b0010011 : word = 9'b1_1111_0010;
						7'b0010001 : word = 9'b1_1111_0011;
						7'b0001111 : word = 9'b1_1111_0100;
						7'b0001101 : word = 9'b1_1111_0101;
						7'b0001011 : word = 9'b1_1111_0110;
						7'b0001001 : word = 9'b1_1111_0111;
						7'b0000111 : word = 9'b1_1111_1000;
						7'b0000110 : word = 9'b1_1111_1001;
						7'b0000100 : word = 9'b1_1111_1010;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd8 : begin
					case (buffer[11:4])
						8'b10010010 : word = 9'b1_0000_0100;
						8'b10000010 : word = 9'b1_0001_0101;
						8'b01111010 : word = 9'b1_0001_0110;
						8'b00101010 : word = 9'b1_0001_1111;
						8'b10000000 : word = 9'b1_0010_0101;
						8'b01111000 : word = 9'b1_0010_0110;
						8'b10000110 : word = 9'b1_0011_0100;
						8'b01111101 : word = 9'b1_0011_0101;
						8'b01110100 : word = 9'b1_0011_0110;
						8'b10010011 : word = 9'b1_0100_0000;
						8'b10000111 : word = 9'b1_0100_0011;
						8'b01111111 : word = 9'b1_0100_0100;
						8'b01110110 : word = 9'b1_0100_0101;
						8'b01110000 : word = 9'b1_0100_0110;
						8'b10000001 : word = 9'b1_0101_0010;
						8'b01111110 : word = 9'b1_0101_0011;
						8'b01110111 : word = 9'b1_0101_0100;
						8'b01110010 : word = 9'b1_0101_0101;
						8'b01111011 : word = 9'b1_0110_0001;
						8'b01111001 : word = 9'b1_0110_0010;
						8'b01110101 : word = 9'b1_0110_0011;
						8'b01110001 : word = 9'b1_0110_0100;
						8'b01110011 : word = 9'b1_0111_0001;
						8'b01101111 : word = 9'b1_0111_0010;
						8'b01101101 : word = 9'b1_0111_0011;
						8'b00010001 : word = 9'b1_0111_1111;
						8'b00010000 : word = 9'b1_1000_1111;
						8'b00001011 : word = 9'b1_1001_1111;
						8'b00001010 : word = 9'b1_1010_1111;
						8'b00000110 : word = 9'b1_1011_1111;
						8'b00000100 : word = 9'b1_1100_1111;
						8'b00000010 : word = 9'b1_1101_1111;
						8'b00000000 : word = 9'b1_1110_1111;
						8'b00101011 : word = 9'b1_1111_0000;
						8'b00000111 : word = 9'b1_1111_1011;
						8'b00000101 : word = 9'b1_1111_1100;
						8'b00000011 : word = 9'b1_1111_1101;
						8'b00000001 : word = 9'b1_1111_1110;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd9 : begin
					case (buffer[11:3])
						9'b100000110 : word = 9'b1_0000_0101;
						9'b011111000 : word = 9'b1_0000_0110;
						9'b001011000 : word = 9'b1_0000_1111;
						9'b011011000 : word = 9'b1_0001_0111;
						9'b011010001 : word = 9'b1_0001_1000;
						9'b011000110 : word = 9'b1_0001_1001;
						9'b011011101 : word = 9'b1_0010_0111;
						9'b011001111 : word = 9'b1_0010_1000;
						9'b011000010 : word = 9'b1_0010_1001;
						9'b010110110 : word = 9'b1_0010_1010;
						9'b011011100 : word = 9'b1_0011_0111;
						9'b011001100 : word = 9'b1_0011_1000;
						9'b010111110 : word = 9'b1_0011_1001;
						9'b010110010 : word = 9'b1_0011_1010;
						9'b011010010 : word = 9'b1_0100_0111;
						9'b011001000 : word = 9'b1_0100_1000;
						9'b010111100 : word = 9'b1_0100_1001;
						9'b100000111 : word = 9'b1_0101_0000;
						9'b011010110 : word = 9'b1_0101_0110;
						9'b011001010 : word = 9'b1_0101_0111;
						9'b011000000 : word = 9'b1_0101_1000;
						9'b010110100 : word = 9'b1_0101_1001;
						9'b011111001 : word = 9'b1_0110_0000;
						9'b011010111 : word = 9'b1_0110_0101;
						9'b011001110 : word = 9'b1_0110_0110;
						9'b011000011 : word = 9'b1_0110_0111;
						9'b010111001 : word = 9'b1_0110_1000;
						9'b011010011 : word = 9'b1_0111_0100;
						9'b011001011 : word = 9'b1_0111_0101;
						9'b011000100 : word = 9'b1_0111_0110;
						9'b010111011 : word = 9'b1_0111_0111;
						9'b011010100 : word = 9'b1_1000_0001;
						9'b011010000 : word = 9'b1_1000_0010;
						9'b011001101 : word = 9'b1_1000_0011;
						9'b011001001 : word = 9'b1_1000_0100;
						9'b011000001 : word = 9'b1_1000_0101;
						9'b010111010 : word = 9'b1_1000_0110;
						9'b010110001 : word = 9'b1_1000_0111;
						9'b010101001 : word = 9'b1_1000_1000;
						9'b011000111 : word = 9'b1_1001_0001;
						9'b011000101 : word = 9'b1_1001_0010;
						9'b010111111 : word = 9'b1_1001_0011;
						9'b010111101 : word = 9'b1_1001_0100;
						9'b010110101 : word = 9'b1_1001_0101;
						9'b010101110 : word = 9'b1_1001_0110;
						9'b010111000 : word = 9'b1_1010_0001;
						9'b010110111 : word = 9'b1_1010_0010;
						9'b010110011 : word = 9'b1_1010_0011;
						9'b010101111 : word = 9'b1_1010_0100;
						9'b010101011 : word = 9'b1_1011_0010;
						9'b010101000 : word = 9'b1_1011_0011;
						9'b010100100 : word = 9'b1_1011_0100;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd10 : begin
					case (buffer[11:2])
						10'b0110110010 : word = 9'b1_0000_0111;
						10'b0110101010 : word = 9'b1_0000_1000;
						10'b0101000111 : word = 9'b1_0001_1010;
						10'b0101011001 : word = 9'b1_0001_1011;
						10'b0100111111 : word = 9'b1_0001_1100;
						10'b0100101001 : word = 9'b1_0001_1101;
						10'b0100010111 : word = 9'b1_0001_1110;
						10'b0101010100 : word = 9'b1_0010_1011;
						10'b0100111011 : word = 9'b1_0010_1100;
						10'b0100100111 : word = 9'b1_0010_1101;
						10'b0101000101 : word = 9'b1_0011_1011;
						10'b0100110111 : word = 9'b1_0011_1100;
						10'b0100100101 : word = 9'b1_0011_1101;
						10'b0100001111 : word = 9'b1_0011_1110;
						10'b0101100000 : word = 9'b1_0100_1010;
						10'b0101000011 : word = 9'b1_0100_1011;
						10'b0100110010 : word = 9'b1_0100_1100;
						10'b0100011101 : word = 9'b1_0100_1101;
						10'b0101010101 : word = 9'b1_0101_1010;
						10'b0100111101 : word = 9'b1_0101_1011;
						10'b0100101101 : word = 9'b1_0101_1100;
						10'b0100011001 : word = 9'b1_0101_1101;
						10'b0100000110 : word = 9'b1_0101_1110;
						10'b0101011011 : word = 9'b1_0110_1001;
						10'b0101001010 : word = 9'b1_0110_1010;
						10'b0100110100 : word = 9'b1_0110_1011;
						10'b0100100011 : word = 9'b1_0110_1100;
						10'b0100010000 : word = 9'b1_0110_1101;
						10'b0110110011 : word = 9'b1_0111_0000;
						10'b0101100001 : word = 9'b1_0111_1000;
						10'b0101001100 : word = 9'b1_0111_1001;
						10'b0100111001 : word = 9'b1_0111_1010;
						10'b0100101010 : word = 9'b1_0111_1011;
						10'b0100011011 : word = 9'b1_0111_1100;
						10'b0110101011 : word = 9'b1_1000_0000;
						10'b0101000000 : word = 9'b1_1000_1001;
						10'b0100101111 : word = 9'b1_1000_1010;
						10'b0100011110 : word = 9'b1_1000_1011;
						10'b0100001100 : word = 9'b1_1000_1100;
						10'b0101001111 : word = 9'b1_1001_0000;
						10'b0101001101 : word = 9'b1_1001_0111;
						10'b0101000001 : word = 9'b1_1001_1000;
						10'b0100110001 : word = 9'b1_1001_1001;
						10'b0100100001 : word = 9'b1_1001_1010;
						10'b0100010011 : word = 9'b1_1001_1011;
						10'b0101011000 : word = 9'b1_1010_0101;
						10'b0101001011 : word = 9'b1_1010_0110;
						10'b0100111010 : word = 9'b1_1010_0111;
						10'b0100110000 : word = 9'b1_1010_1000;
						10'b0100100010 : word = 9'b1_1010_1001;
						10'b0100010101 : word = 9'b1_1010_1010;
						10'b0101011010 : word = 9'b1_1011_0001;
						10'b0100111110 : word = 9'b1_1011_0101;
						10'b0100110101 : word = 9'b1_1011_0110;
						10'b0100101011 : word = 9'b1_1011_0111;
						10'b0100011111 : word = 9'b1_1011_1000;
						10'b0100010100 : word = 9'b1_1011_1001;
						10'b0100000111 : word = 9'b1_1011_1010;
						10'b0101000010 : word = 9'b1_1100_0001;
						10'b0100111100 : word = 9'b1_1100_0010;
						10'b0100111000 : word = 9'b1_1100_0011;
						10'b0100110011 : word = 9'b1_1100_0100;
						10'b0100101110 : word = 9'b1_1100_0101;
						10'b0100100100 : word = 9'b1_1100_0110;
						10'b0100011100 : word = 9'b1_1100_0111;
						10'b0100001101 : word = 9'b1_1100_1000;
						10'b0100000101 : word = 9'b1_1100_1001;
						10'b0100101100 : word = 9'b1_1101_0001;
						10'b0100101000 : word = 9'b1_1101_0010;
						10'b0100100110 : word = 9'b1_1101_0011;
						10'b0100100000 : word = 9'b1_1101_0100;
						10'b0100011010 : word = 9'b1_1101_0101;
						10'b0100010001 : word = 9'b1_1101_0110;
						10'b0100001010 : word = 9'b1_1101_0111;
						10'b0100011000 : word = 9'b1_1110_0001;
						10'b0100010110 : word = 9'b1_1110_0010;
						10'b0100010010 : word = 9'b1_1110_0011;
						10'b0100001011 : word = 9'b1_1110_0100;
						10'b0100001000 : word = 9'b1_1110_0101;
						10'b0100000011 : word = 9'b1_1110_0110;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd11 : begin
					case (buffer[11:1])
						11'b01010011101 : word = 9'b1_0000_1001;
						11'b01010001101 : word = 9'b1_0000_1010;
						11'b01010001001 : word = 9'b1_0000_1011;
						11'b01001101101 : word = 9'b1_0000_1100;
						11'b01000000101 : word = 9'b1_0000_1101;
						11'b01000011101 : word = 9'b1_0010_1110;
						11'b01000011100 : word = 9'b1_0100_1110;
						11'b01000001000 : word = 9'b1_0110_1110;
						11'b01000010011 : word = 9'b1_0111_1101;
						11'b00101111101 : word = 9'b1_0111_1110;
						11'b01000000010 : word = 9'b1_1000_1101;
						11'b00101111001 : word = 9'b1_1000_1110;
						11'b01000001001 : word = 9'b1_1001_1100;
						11'b00101111011 : word = 9'b1_1001_1101;
						11'b00101110011 : word = 9'b1_1001_1110;
						11'b01010011100 : word = 9'b1_1010_0000;
						11'b01000010010 : word = 9'b1_1010_1011;
						11'b00101111111 : word = 9'b1_1010_1100;
						11'b00101110101 : word = 9'b1_1010_1101;
						11'b00101101110 : word = 9'b1_1010_1110;
						11'b01010001100 : word = 9'b1_1011_0000;
						11'b01000000001 : word = 9'b1_1011_1011;
						11'b00101110111 : word = 9'b1_1011_1100;
						11'b00101110000 : word = 9'b1_1011_1101;
						11'b00101101010 : word = 9'b1_1011_1110;
						11'b01010001000 : word = 9'b1_1100_0000;
						11'b01000000000 : word = 9'b1_1100_1010;
						11'b00101111000 : word = 9'b1_1100_1011;
						11'b00101110010 : word = 9'b1_1100_1100;
						11'b00101101100 : word = 9'b1_1100_1101;
						11'b00101100111 : word = 9'b1_1100_1110;
						11'b01001101100 : word = 9'b1_1101_0000;
						11'b01000000011 : word = 9'b1_1101_1000;
						11'b00101111100 : word = 9'b1_1101_1001;
						11'b00101110110 : word = 9'b1_1101_1010;
						11'b00101110001 : word = 9'b1_1101_1011;
						11'b00101101101 : word = 9'b1_1101_1100;
						11'b00101101001 : word = 9'b1_1101_1101;
						11'b00101100101 : word = 9'b1_1101_1110;
						11'b00101111110 : word = 9'b1_1110_0111;
						11'b00101111010 : word = 9'b1_1110_1000;
						11'b00101110100 : word = 9'b1_1110_1001;
						11'b00101101111 : word = 9'b1_1110_1010;
						11'b00101101011 : word = 9'b1_1110_1011;
						11'b00101101000 : word = 9'b1_1110_1100;
						11'b00101100110 : word = 9'b1_1110_1101;
						11'b00101100100 : word = 9'b1_1110_1110;
						default : word = 9'b0_0000_0000;
					endcase
				end
			5'd12 : begin
					case (buffer[11:0])
						12'b010000001000 : word = 9'b1_0000_1110;
						12'b010000001001 : word = 9'b1_1110_0000;
						default : word = 9'b0_0000_0000;
					endcase
				end
			default : word = 9'b0_0000_0000;
		endcase
	end
endmodule


`default_nettype wire
