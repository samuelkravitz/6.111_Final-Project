`default_nettype none
`timescale 1ns / 1ps

module antialias_reorder_tb;

logic clk;
logic rst;

logic window_switching_flag_in;
logic [1:0] block_type_in;
logic mixed_block_flag_in;

logic si_valid;

logic [31:0] ch1_in;
logic [31:0] ch2_in;
logic [9:0] is_pos_in;
logic din_v;

logic [31:0] ch1_x_out, ch1_y_out;
logic [31:0] ch2_x_out, ch2_y_out;
logic [9:0] is_pos_out_x, is_pos_out_y;
logic dout_v;


logic [575:0][31:0] ch1_code, ch2_code;


antialias aliaser_gr1 (
    .clk(clk),
    .rst(rst),
    .window_switching_flag_in(window_switching_flag_in),
    .block_type_in(block_type_in),
    .mixed_block_flag_in(mixed_block_flag_in),
    .new_frame_start(si_valid),
    .ch1_in(ch1_in),
    .ch2_in(ch2_in),
    .din_v(din_v),

    .ch1_out_x(ch1_x_out),
    .ch1_out_y(ch1_y_out),
    .ch2_out_x(ch2_x_out),
    .ch2_out_y(ch2_y_out),

    .is_pos_out_x(is_pos_out_x),
    .is_pos_out_y(is_pos_out_y),
    .dout_v(dout_v)
  );

  antialias aliaser_gr2 (
      .clk(clk),
      .rst(rst),
      .window_switching_flag_in(window_switching_flag_in),
      .block_type_in(block_type_in),
      .mixed_block_flag_in(mixed_block_flag_in),
      .new_frame_start(si_valid),
      .ch1_in(ch1_in),
      .ch2_in(ch2_in),
      .din_v(din_v),

      .ch1_out_x(ch1_x_out),
      .ch1_out_y(ch1_y_out),
      .ch2_out_x(ch2_x_out),
      .ch2_out_y(ch2_y_out),

      .is_pos_out_x(is_pos_out_x),
      .is_pos_out_y(is_pos_out_y),
      .dout_v(dout_v)
    );

logic signed [31:0] ch1_OUT, ch2_OUT;
logic alias_reorder_valid;

antialias_reorder reorderer (
    .clk(clk),
    .rst(rst),
    .ch1_x_in(ch1_x_out),
    .ch1_y_in(ch1_y_out),
    .ch2_x_in(ch2_x_out),
    .ch2_y_in(ch2_y_out),
    .x_pos_in(is_pos_out_x),
    .y_pos_in(is_pos_out_y),
    .valid_in(dout_v),
    .ch1_out(ch1_OUT),
    .ch2_out(ch2_OUT),
    .valid_out(alias_reorder_valid)
  );


granule_assembler UUT (

  );


always begin
  #10;
  clk = !clk;     //clock cycles now happend every 20!
end


initial begin
  $dumpfile("sim/granule_assembler_tb.vcd");
  $dumpvars(0, granule_assembler_tb);
  $display("Starting Sim");

  ch1_code = 18432'h001879cd000e411f00000000fff1bee1ffdc14cbffcfa274ffc2532cffc2532cffc2532cffc2532cffcfa274ffdc14cbffe78633fff1bee1fffa57d9fffa57d9fffa57d9fffa57d9000e411f000e411f0005a8270005a8270005a8270005a827000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f0005a8270005a827fffa57d9fffa57d9000e411f001879cd001879cd001879cd001879cd000e411f000e411f000e411f000e411f0005a8270005a82700000000000000000000000000000000fffa57d9fffa57d9fffa57d9000e411f0005a8270005a82700000000fffa57d9fffa57d9fff1bee1fff1bee1fff1bee1fff1bee1fff1bee1fff1bee1fff1bee1fffa57d9fffa57d9fffa57d9fffa57d9fffa57d9000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f0005a8270005a8270005a8270005a8270005a8270005a8270005a8270005a8270005a8270005a827fffa57d9fffa57d9fffa57d9fffa57d9fffa57d9000000000000000000000000000000000000000000000000000000000005a8270005a8270005a827000e411f000e411f000e411fffe78633ffe78633ffe78633ffe78633fff1bee1fffa57d9fffa57d9000000000005a827000e411f000e411f000e411f000e411f000e411f0005a8270005a82700000000fffa57d9000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f0005a8270005a8270000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  ch2_code = 18432'h001879cd000e411f00000000fff1bee1ffdc14cbffcfa274ffc2532cffc2532cffc2532cffc2532cffcfa274ffdc14cbffe78633fff1bee1fffa57d9fffa57d9fffa57d9fffa57d9000e411f000e411f0005a8270005a8270005a8270005a827000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f0005a8270005a827fffa57d9fffa57d9000e411f001879cd001879cd001879cd001879cd000e411f000e411f000e411f000e411f0005a8270005a82700000000000000000000000000000000fffa57d9fffa57d9fffa57d9000e411f0005a8270005a82700000000fffa57d9fffa57d9fff1bee1fff1bee1fff1bee1fff1bee1fff1bee1fff1bee1fff1bee1fffa57d9fffa57d9fffa57d9fffa57d9fffa57d9000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f0005a8270005a8270005a8270005a8270005a8270005a8270005a8270005a8270005a8270005a827fffa57d9fffa57d9fffa57d9fffa57d9fffa57d9000000000000000000000000000000000000000000000000000000000005a8270005a8270005a827000e411f000e411f000e411fffe78633ffe78633ffe78633ffe78633fff1bee1fffa57d9fffa57d9000000000005a827000e411f000e411f000e411f000e411f000e411f0005a8270005a82700000000fffa57d9000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f000e411f0005a8270005a8270000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

  clk = 0;

  window_switching_flag_in = 1;
  block_type_in = 1;
  mixed_block_flag_in = 0;
  si_valid = 0;

  is_pos_in = 0;
  din_v = 0;

  rst = 0;
  #20;
  rst = 1;
  #20;
  rst = 0;
  #20;

  din_v = 1;
  for (int i = 0; i < 576; i++) begin
    ch1_in = ch1_code[575 - i];
    ch2_in = ch2_code[575 - i];
    is_pos_in = i;
    #20;
  end
  din_v = 0;

  #40000;


  $display("Finishing Sim");
  $finish;

end
endmodule

`default_nettype wire
