`default_nettype none
`timescale 1ns / 1ps



`default_nettype wire
