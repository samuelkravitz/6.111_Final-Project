`default_nettype none
`timescale 1ns / 1ps

module sf_parser_tb;

logic clk;
logic rst;

logic [1037:0] bit_code;
logic [2514:0] bit_code_2;
logic [3202:0] bit_code_3;

logic [1:0][1:0][11:0] part2_3_length;
logic [1:0][1:0][3:0] scalefac_compress;
logic [1:0][1:0]window_switching_flag;
logic [1:0][1:0][1:0] block_type;
logic [1:0][1:0]mixed_block_flag;
logic [1:0][3:0] scfsi;
logic si_valid;

logic [11:0][2:0][3:0] scalefac_s;
logic [20:0][3:0] scalefac_l;
logic axiov;

logic axiid, axiiv;


sf_parser #(.GR(0), .CH(0)) UUT
(
    .clk(clk),
    .rst(rst),
    .axiid(axiid),
    .axiiv(axiiv),

    .scalefac_compress_in(scalefac_compress[0][0]),
    .window_switching_flag_in(window_switching_flag[0][0]),
    .block_type_in(block_type[0][0]),
    .mixed_block_flag_in(mixed_block_flag[0][0]),
    .scfsi_in(scfsi[0]),
    .si_valid(si_valid),
    .scalefac_s(scalefac_s),
    .scalefac_l(scalefac_l),
    .axiov(axiov)
  );

//////////////////////////////////////////

  always begin
    #10;
    clk = !clk;     //clock cycles now happend every 20!
  end

  initial begin
    $dumpfile("sim/sf_parser_sim.vcd");
    $dumpvars(0, sf_parser_tb);
    $display("Starting Sim");

    bit_code_3 = 3203'h002600C940480000424A0100801BCAF31BE88B1E307C1930BF8F8806C419834570B00065A83861001A66885A6271383C5EB0907190E7838A17D494F18392EB8635030C1A1A4250C902329657CAAB9613ABB4672C591940780E1840E4C0518CD50758708422AC530106098B028C98882690291052FF2601891C28998296B80A0C694AA8A5A29D3548359C32558AC99BBAEC46549B72D9BAC201005D52F4F90281644581A8FCFFBF8F55557CBF499034563AEDB9E0236022E9070CAC96248127ED5DB2780A432D999EAB410CBC56A257E0387A36B0101A6BB1771A352DA36FA99762FC8AB139C657946DA64DBC8E1402FDBD142E0C5E56FECA23499680F2804D595DA97B2A6708E0A071AA696C311187A596A59760C8DC0AC8271E79E9981DB85691E2D7DDC745D772E3AFC35F676A08D312B2370E8D1306005E88B0E936662C8F9D97524E5FB74BAC2961BB784FC3F6EC58C7FFFFFFFFE3D3D22BD3D10AEFCB37903B500B7EDFC08ED43B5B3FFFFFFFFF4F82E191035E8283038E38615060A16BB10F920139CB0041C6E24242CC10A504;

    mixed_block_flag = 0;
    scalefac_compress = 16'hffdd;
    window_switching_flag = 4'hf;
    block_type = 8'haa;
    scfsi = 0;

    si_valid = 0;
    axiiv = 0;
    axiid = 0;

    rst = 0;
    clk = 0;
    #20;
    rst = 1;
    #20;
    rst = 0;
    #20;
    si_valid = 1;
    #20;
    si_valid = 0;

    for (int i = 3202; i > 3000; i --) begin
      axiid = bit_code_3[i];
      axiiv = 1;
      #20;
      // axiiv = 0;
      // #80;
    end
    axiiv = 0;
    #2000;

    // bit_code = 1038'b010100100000000000001001100011100110011000100110000111011111000101100001110010111011100111001111011001011000111000011100010010011110000001101010000100100001100101001011011100111000101101001011101000111100111111111011100010000010000001000000010001000001011000010110110011010000000111100000000000010001001000100000000101000011000001011000011010000111100001000001000110001100001001010001100011100001111000101101010010011001101101001010001000000000111101011101100011101000100001010110011000100001000111100010101000101010111011100110001000110110110010011010101110101011011001001010000110101100001001000110100000011100001111001001010000010110001011000101100010101000010111110110101110011011011111101111100010011010101010100001100010101010111001001101010100110111011101111111010010110101001101101010110110001110000111110000111101010111110001011100010001101001000100110100100111101101001111010111000100111101011100010111011101111111110100010011101010111111110111001101011111001111000010010101111001001110010001010010110000100110001101110111001011;
    //
    // gr = 0;
    // mixed_block_flag = 0;
    // scalefac_compress = 5;
    // window_switching_flag = 1;
    // block_type = 3;
    // scfsi = 0;
    // si_valid = 0;
    // axiiv = 0;
    // axiid = 0;
    //
    // rst = 0;
    // clk = 0;
    // #20;
    // rst = 1;
    // #20;
    // rst = 0;
    // #20;
    // si_valid = 1;
    // #20;
    // si_valid = 0;
    // for (int i = 1037; i > 1015; i --) begin
    //   axiid = bit_code[i];
    //   axiiv = 1;
    //   #20;
    //   // axiiv = 0;
    //   // #80;
    // end
    // axiiv = 0;
    // #2000;
    //
    // bit_code_2 = 2515'b0100001000001000001000010111001101100100010101100100010001010110010001001001001011011011001001011101011010111101011001111101010011110110100111010011111101100101110011001001000000110011000001101101000011011001100100000000011000001101000001110100010100100111001100100000011010100000011000001101100110011011001101000000101011010010011001110110010010011011001100000110000110001110000101011010110011100001000011010011010100100011010011000100000010001011100010000001100100110000011101000010011000010000001010001010101010110101000010110011000011000111000011010111101001000000101001011001101010001011110011000010010111011000110101000110100110100110011010000000000100000111101001110101000000100001100101000110011001001110100100001110110110000100101010100101001101110110000011101011101000100001100010001001101110001000000100000011101100010011010110110010100001000000101000101100100011111010110111011101101011011000000110001000010010100111011011100000110101111001000010001101101110100101100010011111010000110000010001000100010100110011000001010000110011100111000001100001010011000011000010111111111011010101010101110111001100010011010000100011100001101010010100001100110100010100101111011111111110101100110011101101100101111011010011110101000111100101001101100000101000000010101101100101000111111101011100010010011001001000011100010000000000010000010101111011110010110001011010100010011100001010010101011010010101100011101001110010011101001010100001010011010001101100110010111011111001010001001000000101100101101101010100010100000110011010000000111111111000111000000101010010001100010101011011000011010010101100111101110000100000101001111001001000101001111010100110111100101110011100101110010011110010001110100010011011100111000101111000000100101100001110101110101100010010000011100110101101101101010001011001110011001101101100000110011110000010001101101110010110110000011101101100011100111010110000011001110000001000011001011100100010000101101100111010011111101110100100011111111010011101101000000111010000011001110111001000111001011111010001010001101110110001010011101100101011100010111011010011001000011000100011000110010110100110100101001101111010110011000110111101000110011001001111101101100001100100000111010001000010011011101001101011110111001001110101010000110001111110101000001101010111001110101100110001101110011011111010010100110101010110011011110000100110101000011100100000000001110110111011100011111111111111110100101101001011100110100110000111111010000101011111001001100011101011000110000000001100100010100001001;
    //
    // gr = 0;
    // mixed_block_flag = 0;
    // scalefac_compress = 15;
    // window_switching_flag = 1;
    // block_type = 2;
    // scfsi = 0;
    // si_valid = 1;
    // axiiv = 0;
    // axiid = 0;
    //
    // for (int i = 2514; i > 2300; i --) begin
    //   axiid = bit_code_2[i];
    //   axiiv = 1;
    //   #20;
    //   if (i==2514) si_valid = 0;
    //   // axiiv = 0;
    //   // #80;
    //
    // end

    $display("Finishing Sim");
    $finish;

  end

endmodule


`default_nettype wire
