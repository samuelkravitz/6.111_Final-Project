`default_nettype none
`timescale 1ns / 1ps

module subband_synth_tb;

logic clk;
logic rst;
logic new_frame_start;
logic [31:0] x_in;
logic x_valid_in;


subband_synthesis UUT (
    clk,
    rst,
    new_frame_start,
    x_in,
    x_valid_in
  );


logic [18431:0] code;

always begin
  #10;
  clk = !clk;     //clock cycles now happend every 20!
end


initial begin
  $dumpfile("sim/subband_synth.vcd");
  $dumpvars(0, subband_synth_tb);
  $display("Starting Sim");

  code = 18432'h00004bf80000ab4f1fffe173000301ce0001a8f01fffff651fffb9391fffbd2200011c5c1fffec9a000572460006f1850000129a1fffbfe11fff676700089cac1fffaeac1fff933f000000691ffffd64000079020003c4881fffeb84000413e21ffff3b61fffb5491fffbf271fffb93c1fff9ea11fffecb60007d5491fffce8b000bf31b000221d61fffec310000096c1fffff861ffffffa1fffc1681fffe5ea1fffca0e1fffeddc1fffb5ef0004a5870003dd011fffbc8b1fff9f1c0007441e00022d84000823bf00052b9a0011a56f000002ce0000adfd1ffffb821ffff2e11ffff7271fffccdd000494231fffecdc0000c19b0000c8af1fffb77a1fffb0db0001058900012fe61fffdb3b000b0dcb1fff5dd01fffd8191fff9c5b1fff993100001c5e0000aec41ffff7b41fffef2d1ffffa900002ac89000012341fffe3cf1fffd6650002d67600024bc51ffffe361fffadd00000d1e8000355a4000256bc1fffad081fffd7631ffffd4b0000bcbc00025ae900018573000255e91ffff8321fffca2e1ffff7711fffd9961fffd6141ffff4d91fffab851ffff1020005a37d0004d32e000a9f8d000599951fffc20f1ffff68d1ffff63600004e821fffe66b000287fa0000b7c9000163de1ffff92a1fffa6050006231b00008e871fffdd161fffe9ef1fff9e3a000512001fffe9dd0004a55c000d86581ffffe931ffff7ee000090ee00009b00000140060000a3401fffe5691fffcd571fffa7801fff9f6b1fffbdfb1fffd6440001399a0003049a0001eb9900028dbd1fffc2b31fffdf601ffffb7e000086e51ffff28900022c661fffbe5100022d9c1fffe62a000076011fffc8300003ce811ffff663000288c71fffbd0d0009e92c1fff91b50003cb921fffbff50006733200000fda0000333100009b5d000092f80001857d0000ec6f00024b400001ab8f000290050002cbeb00022d34000399cc0001c62f0003ac4f0001d2210002bcd0000184d800016b24000028731ffff54f1ffffb0e000148a30002de8b1ffffa591ffff15f1ffff0f5000140c61fffea1f0001399b00016f550000ada61fff912a1fffbedb000164d60005133c1fffc6170000143200005c431ffffb6700000def000220f1000311250001c10500026b9a00059cb000061fdf0003277b0002c0d20005e4400005239b00002c331fffeb460002bccc0001ce9900002df2000054ac1fffecf20002a24c1ffff83d00029f030001e6351fffe1c81fffe7380001b0b0000276181fffd04c1fffaf6f00012bd21fff7a5600055ef51fffd7cd1fffbe3a1ffffedb1fffff6b1ffffbd21ffffa3b1ffffccb1ffff2611ffffca21ffff0261ffff5ba1ffff4c91fffeb581ffffab71fffe5d61ffff8441fffedb51fffed251ffffb991fffe5c800000ac51ffffe6e00003be11ffffb940000704d1ffff84000009d471ffff5460000c4cf1ffff2930000dfa21ffff0910000ee271fffef0e0000e0471fffef1e0000bead1ffff094000019b21ffff97b1ffffaf90000f544000002561fffec14000093c000017f2b1fffea931fffe89e0001f35b0000e7ec1fffd9bb000005a5000309e21fffe9561fffce8000024c9a000024a70000531c1fffed99000072d31fffd5f10001b0ff00009e190001116100026a021fffd5d91fffe9bb1ffff07d1fffcc03000658861fffe93d00052ffe1fffd88b1fffcb870000225c0000b12c000001e9000194bb1ffff903000195d81ffff8480000d5a71fffff771fffff6b000116701ffff3e300030b9f1fffef22000503a60000089f000541c80003130a1fffffb8000012e20001a7060000090f1ffff5bd0003909d0001370d1ffff1450000c7991ffff262000133171fffe17c1fff926e00018c551ffffe341fff88bd1ffff7090000660b1ffffd291fffffd4000031d61fffecaa00005c5f1ffff9e31fffe32e0000e38b1fffe7b31fffe57b0001288a1fffd2c31ffff4410000df011fffc2ad0000e0d01ffffeb41fffbf011ffffe621ffff9d6000046510000f9a7000007771fffeac91ffff7c10001844400013c1a1fffea701fffe0600000cf1700028bfa1ffffedf1fffce831fffec2d0002ecb000024f890000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ffffebe000039091ffff9bd000094a51ffff41f0000d2951ffff31f0000bb061ffff5110000bedd1ffff0c40001436f1fffe6b70001cad61fffe2880001c3bf1fffe4ec0001cc5d00000f451ffff9670000bb241ffff5c3000008120000d77f1fffe81c000178e51ffff5bc1ffff4cc0001eb2d1fffda8000019df80000137e1fffdf8800034c261fffcde500015dc4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

  clk = 0;

  clk = 0;
  rst = 0;
  x_in = 0;
  x_valid_in = 0;
  new_frame_start = 0;

  #20;
  rst = 1;
  #20;
  rst = 0;
  #20;

  x_valid_in = 1;
  for (int i = 0; i < 576; i++) begin
    x_in = code[(18431 - (32 * i))-: 32];
    #20;
  end
  x_valid_in = 0;


  code = 18432'h1fff7b010005b83500020aa01fffa3de1fff7a6f1ffee5601fff8ca00001090700e7b38a00c8b2651fd74a8a1f8bec1e1eedcbbc1ec86f451ed3d36e1f17b03a1f79673c1f9f6b8500002fdd1fffb0611fffd7e4000d027c1ffe859e000935f800017124002785231fff778300d4cf0000ffbaa100e673da005f5c551ff3c1f9012922ea0048ab0c1ff7d0fe010b68b61fffb7580003befe0012905a000bc3040004f509000657cc1fff1c2b1ffdfdf81ffc11171ff537eb1ffb84910114b1e8014018570015b8de1ff2ead71ff81c941ff86f071fffc8851fffd3650007f3d71fffdf1e1fffb80b1ffee77e1fffdebd0008c4201fffe61c003e9d8b000141ac1fefa5c1020f89c81ff691fb1ffaf31c006149ff1feec2cb001451181ffab40c0003944c000739381fffcb171fff796c1ffffb38001094de1fffd23d0009a84d1ffed98b1ff402971ffc2907000be302009d43cb006008251ffa92910040027e1ffe40cf008fab1f000061301fffd7ee1ffff6620009ebb91fffb7731fff52011fff30f11fff2a2d1ff9e53f1ff51720004a87361ff9c7a400168e031ffb4cd20064c3c10064e8b61ffc94481ff6b00e1fffaa471fff5ec81fff16d01fffee991fffdef71fffa3980016756b000906de0058109300146db701caaf941ffb6b6e1ffc314d1ffdda991fff81701ffea8f00048332d005610081fff91471ffffcf91fffe2b20008a8bc0002b0890004d40e1ffe8cf90024c5191ffc814600afd3f000c93b041ff9974200f8c5fe1ff81abf00112d2500369e04007e24a70006617b1fffbc4b1fffb3180008fd6e1fff80c11fffedfc1fff7dbe000484d8000541ef0006d4731ffb309b1ffd5a9a007b365100159c841ffe18a01ffe3a69005766a50028c19a1ffff21600002d3200010ed01fffd13200014f1a1fff7d710002003a0000b9b21fffd75e1ffee9021fffa8251ffec09700626b901fff81331ffdcee0000b2003003572df00b168b21ffec7f81fff98a81fffbcab1ffff83b1fffbfc3000153430007222b1fffc82100069273003374591ffa246d1ff603540056f9541ffef9050131fe92002e9a570069fa9e1ffd13941ffa85c21fffbded1fffafbb00026b240003cb7a1fffa83c1fffd27f000a7e25000aedbf1ffe85e60036e42d1ffdd3a70013c1071ffa63fe0012ce931ffc4d8c1ff97b4400906dd2000f42871fff6f0f000463780005970a1fffb4f9000061361ffff2620001f9d600065d7700124643001478cf006a7d6a1ff57d711ffbfaf71ffb110a1fff124f0005b3101ffd7afc1ffe36ed00001ad51fffec7a1ffff7141ffffda81fffe34e1fffda9f1fffa2920004e2401ffbce40000a3aad003ead561fffe306003539fd00094b0d1ffddcfa1ff97b960047c54b001dfdce000091181ffff31e000084481ffff7ad0001d6ad1ffff7bb000b63ec1fffc3160030c1b60033e2b61ffec6371fff9e251ff452f7001cee680043328b1ffec2ea1ff9eeee00287de0000309181fffc1071fffe5e30005fccb1fffeef61fff8a500000f6ff000443721ffe8d560031cfaf1ffc90180001ac6d003b64601ffe1c741ff86a391fffe6631ffec4441ffd7a111fffc0b50000b4191fffde9f000ec0e81fffa45b0009641f1fff0d2a1ffec386000b42fd002797921ffe07ac1fffe7090019754c1ffb86f90024a8ee1fff99180024cef5004bff61000331ce0006be6900004f110008f4be1fffdb8c0009e09c1fffe9d11fffbf0c0009927a001d10ee1ffd95d200232c2d1fffef69000192130034d3471ffee1e31ffdedab1fff97bf00018d6b0003609f1fffb5400009a3fc001122571fff78340008b00c1fffbd41000607dc1fff2be2005a387f1fff1e711fff9fe2001a2a651ffef3d11ffd1013000626e00002f5870002eb2d1fffe1191fffca240005395b1fff9a9d1fffce9f00025ed71ffe7cad1ffdd172000ca11d00287a1d1fff48811ffdd8f9002b399500192bf00013eee50009e7830001dd611fffd25b1fffbd310001b5b000062b790000c4be1fff8c651fffd641000cb30700108a21003ab70d0021c4dc000f86941ffed6ea1fff793d1ffdeb0c1ffeeb911fff7d33001c7713000000000000000000000000000000000000000000000000000324d61ffedbee000f774e001427dd1ffd3ee10017e15d0000d756000098f71ffde3020016594d1ffe47051fffc4b11fffdc820002fc4a1fffc0420004f6e81fffa63a0005a1961fffd41b00092005001431a71ffe3c371fff295a1ffefa46001f3caa1fffc6c21ffe627f1ffed8821fff9d4f1fff122200016c1a1fffbe33000570f41fffb8ff0000cdf60004e8821fff98a1000d6c5c1fffe84a001f7b791fff3cff0026633a1fff4bb20010f8761fff853b1fff4587000257d81ffeff10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

  x_valid_in = 1;
  for (int i = 0; i < 576; i++) begin
    x_in = code[(18431 - (32 * i))-: 32];
    #20;
  end
  x_valid_in = 0;


  #400000;


  $display("Finishing Sim");
  $finish;

end
endmodule

`default_nettype wire
